input wire c1_sys_clk_p;
input wire c1_sys_clk_n;

output c1_ddr4_act_n;
output [16:0] c1_ddr4_adr;
output [1:0] c1_ddr4_ba;
output [0:0] c1_ddr4_bg;
output [0:0] c1_ddr4_cke;
output [0:0] c1_ddr4_odt;
output [0:0] c1_ddr4_cs_n;
output [0:0] c1_ddr4_ck_t;
output [0:0] c1_ddr4_ck_c;
output c1_ddr4_reset_n;
inout [3:0] c1_ddr4_dm_dbi_n;
inout [31:0] c1_ddr4_dq;
inout [3:0] c1_ddr4_dqs_c;
inout [3:0] c1_ddr4_dqs_t;
