	,.ddr3_dq(ddr3_dq)
	,.ddr3_dqs_n(ddr3_dqs_n)
	,.ddr3_dqs_p(ddr3_dqs_p)
	,.ddr3_addr(ddr3_addr)
	,.ddr3_ba(ddr3_ba)
	,.ddr3_ras_n(ddr3_ras_n)
	,.ddr3_cas_n(ddr3_cas_n)
	,.ddr3_we_n(ddr3_we_n)
	,.ddr3_reset_n(ddr3_reset_n)
	,.ddr3_ck_p(ddr3_ck_p)
	,.ddr3_ck_n(ddr3_ck_n)
	,.ddr3_cke(ddr3_cke)
	,.ddr3_cs_n(ddr3_cs_n)
	,.ddr3_dm(ddr3_dm)
	,.ddr3_odt(ddr3_odt)