,.c2_sys_clk_p(c2_sys_clk_p)
,.c2_sys_clk_n(c2_sys_clk_n)

,.c2_ddr3_addr(c2_ddr3_addr)
,.c2_ddr3_ba(c2_ddr3_ba)
,.c2_ddr3_ras_n(c2_ddr3_ras_n)
,.c2_ddr3_cas_n(c2_ddr3_cas_n)
,.c2_ddr3_we_n(c2_ddr3_we_n)
,.c2_ddr3_cke(c2_ddr3_cke)
,.c2_ddr3_odt(c2_ddr3_odt)
,.c2_ddr3_cs_n(c2_ddr3_cs_n)
,.ddrx_rtl_0_ck_p(ddrx_rtl_0_ck_p)
,.ddrx_rtl_0_ck_n(ddrx_rtl_0_ck_n)
,.c2_ddr3_reset_n(c2_ddr3_reset_n)
,.c2_ddr3_dm(c2_ddr3_dm)
,.c2_ddr3_dq(c2_ddr3_dq)
,.c2_ddr3_dqs_p(c2_ddr3_dqs_p)
,.c2_ddr3_dqs_n(c2_ddr3_dqs_n)
