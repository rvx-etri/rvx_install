input wire c2_sys_clk_p;
input wire c2_sys_clk_n;

output wire [14:0] c2_ddr3_addr;
output wire [2:0] c2_ddr3_ba;
output wire c2_ddr3_ras_n;
output wire c2_ddr3_cas_n;
output wire c2_ddr3_we_n;
output wire [0:0] c2_ddr3_cke;
output wire [0:0] c2_ddr3_odt;
output wire [0:0] c2_ddr3_cs_n;
output wire [0:0] ddrx_rtl_0_ck_p;
output wire [0:0] ddrx_rtl_0_ck_n;
output wire c2_ddr3_reset_n;
output wire [3:0] c2_ddr3_dm;
inout wire [31:0] c2_ddr3_dq;
inout wire [3:0] c2_ddr3_dqs_p;
inout wire [3:0] c2_ddr3_dqs_n;
