,.c1_sys_clk_p(c1_sys_clk_p)
,.c1_sys_clk_n(c1_sys_clk_n)

,.c1_ddr4_act_n(c1_ddr4_act_n)
,.c1_ddr4_adr(c1_ddr4_adr)
,.c1_ddr4_ba(c1_ddr4_ba)
,.c1_ddr4_bg(c1_ddr4_bg)
,.c1_ddr4_cke(c1_ddr4_cke)
,.c1_ddr4_odt(c1_ddr4_odt)
,.c1_ddr4_cs_n(c1_ddr4_cs_n)
,.c1_ddr4_ck_t(c1_ddr4_ck_t)
,.c1_ddr4_ck_c(c1_ddr4_ck_c)
,.c1_ddr4_reset_n(c1_ddr4_reset_n)
,.c1_ddr4_dm_dbi_n(c1_ddr4_dm_dbi_n)
,.c1_ddr4_dq(c1_ddr4_dq)
,.c1_ddr4_dqs_c(c1_ddr4_dqs_c)
,.c1_ddr4_dqs_t(c1_ddr4_dqs_t)
